library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

entity Picture_Block_RAM is
	generic (
		AddressWidth : integer := 16;
		DataWidth : integer := 12
	);
	port (
		CLK : in std_logic;
		WR : in std_logic;
		AB : in std_logic_vector(AddressWidth - 1 downto 0);
		DB : out std_logic_vector(DataWidth - 1 downto 0)
	);
end Picture_Block_RAM;	

architecture Behavioral of Picture_Block_RAM is

	subtype word is std_logic_vector (DataWidth - 1 downto 0);
	
	type tram is array (0 to 3599) of word;
	
	constant picture : tram := (
	"011001011110",
"101110111101",
"101010101101",
"110111011101",
"110111011101",
"101010101101",
"101110101101",
"011001101110",
"010101011101",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"010001001100",
"011001101111",
"101110111111",
"011101111111",
"111011101111",
"111011011111",
"011101111111",
"101110111111",
"011101111111",
"010000111111",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"011001101111",
"100110011111",
"011101111111",
"110011001111",
"101110111111",
"100001111111",
"100110011111",
"011101111111",
"010000111110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"011001101111",
"011101111111",
"110011001111",
"101010011111",
"101010011111",
"110011001111",
"011101111111",
"011101111111",
"010000111110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"010101011110",
"100010001111",
"111111111111",
"100010001111",
"100110011111",
"111111111111",
"011101111111",
"011001101111",
"010000111110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"010101011110",
"100110011111",
"111111111111",
"100010001111",
"100110011111",
"111111111111",
"100010001111",
"011001101111",
"010000111110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"010101011110",
"011101111111",
"111011101111",
"100010001111",
"100110011111",
"111011101111",
"011101101111",
"011001101111",
"010000111110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"011001101111",
"100010001111",
"101010101111",
"101010101111",
"101010101111",
"101110101111",
"100010001111",
"011101111111",
"010000111110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"011001101111",
"101010101111",
"011001101111",
"110111011111",
"110011001111",
"011101101111",
"101010101111",
"011101111111",
"010000111110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"011001101111",
"110011001111",
"100010001111",
"111111111111",
"111011101111",
"100010001111",
"110011001111",
"011101111111",
"010000111110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"011001101111",
"101010101111",
"110011001111",
"110111011111",
"110111011111",
"110011001111",
"101010101111",
"011101111111",
"010000111110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"011001011111",
"010101011111",
"100010001111",
"100010001111",
"100010001111",
"100110001111",
"010101011111",
"011101101111",
"010000111110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"010101011110",
"010101001111",
"010101011111",
"011101101111",
"011001101111",
"011001011111",
"010001001111",
"011001101111",
"010000111110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"011001011111",
"010101011111",
"100010001111",
"100010001111",
"100010001111",
"100110011111",
"010101011111",
"011101101111",
"010000111110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"011001101111",
"101010101111",
"111011101111",
"110111011111",
"110111011111",
"111011101111",
"101010101111",
"011101111111",
"010000111110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"011001101111",
"110111011111",
"111111111111",
"111111111111",
"111111111111",
"111111111111",
"110011001111",
"011101111111",
"010000111110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"011001101111",
"110011001111",
"110011001111",
"111111111111",
"111111111111",
"110011001111",
"110011001111",
"011101111111",
"010000111110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"011001101111",
"110011001111",
"011101101111",
"111011101111",
"111011101111",
"011101101111",
"101110111111",
"011101111111",
"010000111110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"011001101111",
"101010101111",
"001100111110",
"110010111111",
"110011001111",
"001100111110",
"100110001111",
"011101111111",
"010000111110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"011001101111",
"011101111111",
"001000011110",
"100010001111",
"101010011111",
"001000011110",
"011001011111",
"011101111111",
"010000111110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"011001101111",
"011001101111",
"001000011110",
"011101111111",
"100010001111",
"001000011110",
"010001001111",
"011101111111",
"010000111110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"011001101111",
"100110011111",
"100110011111",
"101010011111",
"101010101111",
"100110011111",
"100010001111",
"011101111111",
"010000111110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"011001101111",
"110011001111",
"111111111111",
"101010101111",
"101110111111",
"111111111111",
"110011001111",
"011101111111",
"010000111110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"011001101111",
"110111011111",
"111111111111",
"100010001111",
"100110011111",
"111111111111",
"110011001111",
"011101111111",
"010000111110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"011001101111",
"110111011111",
"111111111111",
"100110011111",
"100110011111",
"111111111111",
"110011001111",
"011101111111",
"010000111110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"011001101111",
"110111011111",
"110111011111",
"101110111111",
"101010101111",
"111011101111",
"110011001111",
"011101111111",
"010000111110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"011001101111",
"110111011111",
"101110111111",
"110111011111",
"110011001111",
"110011001111",
"110111001111",
"011101111111",
"010000111110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"010101011111",
"101110111111",
"101010101111",
"110011001111",
"101110111111",
"101010101111",
"101110111111",
"011001101111",
"010000111110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"010101011110",
"100001111111",
"100110011111",
"100110011111",
"100010001111",
"100110011111",
"011101111111",
"011001101111",
"010000111110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"011001101110",
"010101011111",
"101010101111",
"100110011111",
"100110011111",
"100110011111",
"011001011111",
"011101111111",
"010000111110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"011001101111",
"010101011111",
"101110111111",
"101110111111",
"101110111111",
"101010101111",
"011001101111",
"011101111111",
"010000111110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"011001011111",
"010101011111",
"101010101111",
"100110011111",
"100110011111",
"100110011111",
"011001101111",
"011101111111",
"010000111110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"010101011110",
"100001111111",
"100110011111",
"100110001111",
"100010001111",
"100110011111",
"011001101111",
"011001101111",
"010000111110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"010101011111",
"101110111111",
"101010101111",
"110011001111",
"101110111111",
"101010101111",
"101010101111",
"011001101111",
"010000111110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"011001101111",
"110111011111",
"110011001111",
"110011001111",
"110011001111",
"110011001111",
"110011001111",
"011101111111",
"010000111110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"011001101111",
"110111011111",
"110111011111",
"101010101111",
"101010101111",
"111011101111",
"110011001111",
"011101111111",
"010000111110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"011001101111",
"110111011111",
"111111111111",
"100110001111",
"100110011111",
"111111111111",
"110011001111",
"011101111111",
"010000111110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"011001101111",
"110111011111",
"111111111111",
"100110001111",
"100110011111",
"111111111111",
"110011001111",
"011101111111",
"010000111110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"001000011110",
"011001101111",
"110011001111",
"111111111111",
"101110111111",
"101110111111",
"111111111111",
"110010111111",
"011101111111",
"010000111111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"001000011111",
"011001101111",
"100110001111",
"100010001111",
"101010011111",
"101010101111",
"100010001111",
"011101111111",
"011101111110",
"010101111001",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"001101100111",
"011001101111",
"011001101111",
"000100011110",
"011101111111",
"100010001111",
"000100011110",
"010001001111",
"011101111110",
"011010100011",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"011001101111",
"011101111111",
"001000011110",
"100110001111",
"101010101111",
"001000011110",
"011001101111",
"011101111110",
"011010100011",
"010010100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"011001101111",
"101010101111",
"001100111110",
"110011001111",
"110111011111",
"001100111111",
"100110011111",
"011101111110",
"011010100011",
"010010100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"011001101111",
"110011001111",
"011101111111",
"111011101111",
"111111111111",
"011101111111",
"101110111111",
"011101111110",
"011010100011",
"010010100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"011001101111",
"110011001111",
"110111011111",
"111111111111",
"111111111111",
"110111011111",
"110011001111",
"011101111110",
"011010100011",
"010010100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"011001101111",
"110011001111",
"111111111111",
"111111111111",
"111111111111",
"111111111111",
"110011001111",
"011101111110",
"011010100011",
"010010100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"011001101111",
"100110001111",
"110011001111",
"110011001111",
"110011001111",
"110011001111",
"100010001111",
"011101111110",
"011010100011",
"010010100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010101011110",
"010001001111",
"011101111111",
"100001111111",
"011101111111",
"011101111111",
"010001001111",
"011101111110",
"011010100011",
"010010100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010101011110",
"010101001111",
"011001011111",
"011101101111",
"011001101111",
"011001101111",
"010001001111",
"011001101110",
"011010100011",
"010010100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"011001101111",
"011001101111",
"101010101111",
"101010101111",
"100110011111",
"101010101111",
"011001101111",
"011101111110",
"011010100011",
"010010100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"011001101111",
"101110111111",
"110011001111",
"111011101111",
"111011101111",
"110011001111",
"101110111111",
"011101111110",
"011010100011",
"010010100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"011001101111",
"101110111111",
"011101101111",
"111011101111",
"111011101111",
"011101111111",
"101110111111",
"011101111110",
"011010100011",
"010010100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"011001101111",
"100110011111",
"011101111111",
"110011001111",
"110010111111",
"011101111111",
"100110011111",
"011101111110",
"011010100011",
"010010100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"011001101111",
"011101111111",
"110011001111",
"101010101111",
"101010101111",
"110011001111",
"011101111111",
"011101111110",
"011010100011",
"010010100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010101011110",
"011101111111",
"111111111111",
"100010001111",
"100110011111",
"111111111111",
"011101111111",
"011001101110",
"011010100011",
"010010100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010101011110",
"100110011111",
"111111111111",
"100010001111",
"100110011111",
"111111111111",
"100010001111",
"011001101110",
"011010100011",
"010010100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010101011110",
"011101111111",
"111011101111",
"100010001111",
"100110011111",
"111011101111",
"011101101111",
"011001111110",
"011010100011",
"010010100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"011001101111",
"100001111111",
"101110111111",
"101010101111",
"101010101111",
"101110111111",
"011101111111",
"011101111110",
"011010100011",
"010010100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"011001101111",
"101010101111",
"011101101111",
"110111011111",
"110011001111",
"011101101111",
"101010101111",
"011101111110",
"011010100011",
"010010100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"011001101111",
"110011001111",
"011101111111",
"111011101111",
"111011101111",
"100001111111",
"110010111111",
"011101111110",
"011010100011",
"010010100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000",
"010110100000"
	);	
	
	signal adrreg : natural;
	signal rom_data : std_logic_vector(DataWidth - 1 downto 0);
	signal reg_out : std_logic_vector(DataWidth - 1 downto 0);

begin
	
	adrreg <= to_integer(unsigned(AB));
	rom_data <= picture(adrreg);
	
	P_REG_OUT: process (CLK,WR,rom_data)
	begin
		if (WR= '1') then
			if (rising_edge (CLK)) then
				reg_out<=rom_data;
			end if;
		end if;
	end process;
	
	DB <= reg_out;
end Behavioral;

